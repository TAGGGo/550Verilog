module left_shift(opA, amt, cout);
	input [31:0] opA;
	input [4:0] amt;
	output [31:0] cout;
	wire zero;
	assign zero = 1'b0;
	
	// if amt == 0, choose lower indexed bit
	
	// layer 1
	wire [31:0] tmp_1;
	my_mux my_mux1(opA[31], opA[30], amt[0], tmp_1[31]);
	my_mux my_mux2(opA[30], opA[29], amt[0], tmp_1[30]);
	my_mux my_mux3(opA[29], opA[28], amt[0], tmp_1[29]);
	my_mux my_mux4(opA[28], opA[27], amt[0], tmp_1[28]);
	my_mux my_mux5(opA[27], opA[26], amt[0], tmp_1[27]);
	my_mux my_mux6(opA[26], opA[25], amt[0], tmp_1[26]);
	my_mux my_mux7(opA[25], opA[24], amt[0], tmp_1[25]);
	my_mux my_mux8(opA[24], opA[23], amt[0], tmp_1[24]);
	my_mux my_mux9(opA[23], opA[22], amt[0], tmp_1[23]);
	my_mux my_mux10(opA[22], opA[21], amt[0], tmp_1[22]);
	my_mux my_mux11(opA[21], opA[20], amt[0], tmp_1[21]);
	my_mux my_mux12(opA[20], opA[19], amt[0], tmp_1[20]);
	my_mux my_mux13(opA[19], opA[18], amt[0], tmp_1[19]);
	my_mux my_mux14(opA[18], opA[17], amt[0], tmp_1[18]);
	my_mux my_mux15(opA[17], opA[16], amt[0], tmp_1[17]);
	my_mux my_mux16(opA[16], opA[15], amt[0], tmp_1[16]);
	my_mux my_mux17(opA[15], opA[14], amt[0], tmp_1[15]);
	my_mux my_mux18(opA[14], opA[13], amt[0], tmp_1[14]);
	my_mux my_mux19(opA[13], opA[12], amt[0], tmp_1[13]);
	my_mux my_mux20(opA[12], opA[11], amt[0], tmp_1[12]);
	my_mux my_mux21(opA[11], opA[10], amt[0], tmp_1[11]);
	my_mux my_mux22(opA[10], opA[9], amt[0], tmp_1[10]);
	my_mux my_mux23(opA[9], opA[8], amt[0], tmp_1[9]);
	my_mux my_mux24(opA[8], opA[7], amt[0], tmp_1[8]);
	my_mux my_mux25(opA[7], opA[6], amt[0], tmp_1[7]);
	my_mux my_mux26(opA[6], opA[5], amt[0], tmp_1[6]);
	my_mux my_mux27(opA[5], opA[4], amt[0], tmp_1[5]);
	my_mux my_mux28(opA[4], opA[3], amt[0], tmp_1[4]);
	my_mux my_mux29(opA[3], opA[2], amt[0], tmp_1[3]);
	my_mux my_mux30(opA[2], opA[1], amt[0], tmp_1[2]);
	my_mux my_mux31(opA[1], opA[0], amt[0], tmp_1[1]);
	my_mux my_mux32(opA[0], zero, amt[0], tmp_1[0]);
	
	// layer 2
	wire [31:0] tmp_2;
	my_mux my_mux33(tmp_1[31], tmp_1[29], amt[1], tmp_2[31]);
	my_mux my_mux34(tmp_1[30], tmp_1[28], amt[1], tmp_2[30]);
	my_mux my_mux35(tmp_1[29], tmp_1[27], amt[1], tmp_2[29]);
	my_mux my_mux36(tmp_1[28], tmp_1[26], amt[1], tmp_2[28]);
	my_mux my_mux37(tmp_1[27], tmp_1[25], amt[1], tmp_2[27]);
	my_mux my_mux38(tmp_1[26], tmp_1[24], amt[1], tmp_2[26]);
	my_mux my_mux39(tmp_1[25], tmp_1[23], amt[1], tmp_2[25]);
	my_mux my_mux40(tmp_1[24], tmp_1[22], amt[1], tmp_2[24]);
	my_mux my_mux41(tmp_1[23], tmp_1[21], amt[1], tmp_2[23]);
	my_mux my_mux42(tmp_1[22], tmp_1[20], amt[1], tmp_2[22]);
	my_mux my_mux43(tmp_1[21], tmp_1[19], amt[1], tmp_2[21]);
	my_mux my_mux44(tmp_1[20], tmp_1[18], amt[1], tmp_2[20]);
	my_mux my_mux45(tmp_1[19], tmp_1[17], amt[1], tmp_2[19]);
	my_mux my_mux46(tmp_1[18], tmp_1[16], amt[1], tmp_2[18]);
	my_mux my_mux47(tmp_1[17], tmp_1[15], amt[1], tmp_2[17]);
	my_mux my_mux48(tmp_1[16], tmp_1[14], amt[1], tmp_2[16]);
	my_mux my_mux49(tmp_1[15], tmp_1[13], amt[1], tmp_2[15]);
	my_mux my_mux50(tmp_1[14], tmp_1[12], amt[1], tmp_2[14]);
	my_mux my_mux51(tmp_1[13], tmp_1[11], amt[1], tmp_2[13]);
	my_mux my_mux52(tmp_1[12], tmp_1[10], amt[1], tmp_2[12]);
	my_mux my_mux53(tmp_1[11], tmp_1[9], amt[1], tmp_2[11]);
	my_mux my_mux54(tmp_1[10], tmp_1[8], amt[1], tmp_2[10]);
	my_mux my_mux55(tmp_1[9], tmp_1[7], amt[1], tmp_2[9]);
	my_mux my_mux56(tmp_1[8], tmp_1[6], amt[1], tmp_2[8]);
	my_mux my_mux57(tmp_1[7], tmp_1[5], amt[1], tmp_2[7]);
	my_mux my_mux58(tmp_1[6], tmp_1[4], amt[1], tmp_2[6]);
	my_mux my_mux59(tmp_1[5], tmp_1[3], amt[1], tmp_2[5]);
	my_mux my_mux60(tmp_1[4], tmp_1[2], amt[1], tmp_2[4]);
	my_mux my_mux61(tmp_1[3], tmp_1[1], amt[1], tmp_2[3]);
	my_mux my_mux62(tmp_1[2], tmp_1[0], amt[1], tmp_2[2]);
	my_mux my_mux63(tmp_1[1], zero, amt[1], tmp_2[1]);
	my_mux my_mux64(tmp_1[0], zero, amt[1], tmp_2[0]);
	
	// layer 3
	wire [31:0] tmp_3;
	my_mux my_mux65(tmp_2[31], tmp_2[27], amt[2], tmp_3[31]);
	my_mux my_mux66(tmp_2[30], tmp_2[26], amt[2], tmp_3[30]);
	my_mux my_mux67(tmp_2[29], tmp_2[25], amt[2], tmp_3[29]);
	my_mux my_mux68(tmp_2[28], tmp_2[24], amt[2], tmp_3[28]);
	my_mux my_mux69(tmp_2[27], tmp_2[23], amt[2], tmp_3[27]);
	my_mux my_mux70(tmp_2[26], tmp_2[22], amt[2], tmp_3[26]);
	my_mux my_mux71(tmp_2[25], tmp_2[21], amt[2], tmp_3[25]);
	my_mux my_mux72(tmp_2[24], tmp_2[20], amt[2], tmp_3[24]);
	my_mux my_mux73(tmp_2[23], tmp_2[19], amt[2], tmp_3[23]);
	my_mux my_mux74(tmp_2[22], tmp_2[18], amt[2], tmp_3[22]);
	my_mux my_mux75(tmp_2[21], tmp_2[17], amt[2], tmp_3[21]);
	my_mux my_mux76(tmp_2[20], tmp_2[16], amt[2], tmp_3[20]);
	my_mux my_mux77(tmp_2[19], tmp_2[15], amt[2], tmp_3[19]);
	my_mux my_mux78(tmp_2[18], tmp_2[14], amt[2], tmp_3[18]);
	my_mux my_mux79(tmp_2[17], tmp_2[13], amt[2], tmp_3[17]);
	my_mux my_mux80(tmp_2[16], tmp_2[12], amt[2], tmp_3[16]);
	my_mux my_mux81(tmp_2[15], tmp_2[11], amt[2], tmp_3[15]);
	my_mux my_mux82(tmp_2[14], tmp_2[10], amt[2], tmp_3[14]);
	my_mux my_mux83(tmp_2[13], tmp_2[9], amt[2], tmp_3[13]);
	my_mux my_mux84(tmp_2[12], tmp_2[8], amt[2], tmp_3[12]);
	my_mux my_mux85(tmp_2[11], tmp_2[7], amt[2], tmp_3[11]);
	my_mux my_mux86(tmp_2[10], tmp_2[6], amt[2], tmp_3[10]);
	my_mux my_mux87(tmp_2[9], tmp_2[5], amt[2], tmp_3[9]);
	my_mux my_mux88(tmp_2[8], tmp_2[4], amt[2], tmp_3[8]);
	my_mux my_mux89(tmp_2[7], tmp_2[3], amt[2], tmp_3[7]);
	my_mux my_mux90(tmp_2[6], tmp_2[2], amt[2], tmp_3[6]);
	my_mux my_mux91(tmp_2[5], tmp_2[1], amt[2], tmp_3[5]);
	my_mux my_mux92(tmp_2[4], tmp_2[0], amt[2], tmp_3[4]);
	my_mux my_mux93(tmp_2[3], zero, amt[2], tmp_3[3]);
	my_mux my_mux94(tmp_2[2], zero, amt[2], tmp_3[2]);
	my_mux my_mux95(tmp_2[1], zero, amt[2], tmp_3[1]);
	my_mux my_mux96(tmp_2[0], zero, amt[2], tmp_3[0]);
	
	// layer 4
	wire [31:0] tmp_4;
	my_mux my_mux97(tmp_3[31], tmp_3[23], amt[3], tmp_4[31]);
	my_mux my_mux98(tmp_3[30], tmp_3[22], amt[3], tmp_4[30]);
	my_mux my_mux99(tmp_3[29], tmp_3[21], amt[3], tmp_4[29]);
	my_mux my_mux100(tmp_3[28], tmp_3[20], amt[3], tmp_4[28]);
	my_mux my_mux101(tmp_3[27], tmp_3[19], amt[3], tmp_4[27]);
	my_mux my_mux102(tmp_3[26], tmp_3[18], amt[3], tmp_4[26]);
	my_mux my_mux103(tmp_3[25], tmp_3[17], amt[3], tmp_4[25]);
	my_mux my_mux104(tmp_3[24], tmp_3[16], amt[3], tmp_4[24]);
	my_mux my_mux105(tmp_3[23], tmp_3[15], amt[3], tmp_4[23]);
	my_mux my_mux106(tmp_3[22], tmp_3[14], amt[3], tmp_4[22]);
	my_mux my_mux107(tmp_3[21], tmp_3[13], amt[3], tmp_4[21]);
	my_mux my_mux108(tmp_3[20], tmp_3[12], amt[3], tmp_4[20]);
	my_mux my_mux109(tmp_3[19], tmp_3[11], amt[3], tmp_4[19]);
	my_mux my_mux110(tmp_3[18], tmp_3[10], amt[3], tmp_4[18]);
	my_mux my_mux111(tmp_3[17], tmp_3[9], amt[3], tmp_4[17]);
	my_mux my_mux112(tmp_3[16], tmp_3[8], amt[3], tmp_4[16]);
	my_mux my_mux113(tmp_3[15], tmp_3[7], amt[3], tmp_4[15]);
	my_mux my_mux114(tmp_3[14], tmp_3[6], amt[3], tmp_4[14]);
	my_mux my_mux115(tmp_3[13], tmp_3[5], amt[3], tmp_4[13]);
	my_mux my_mux116(tmp_3[12], tmp_3[4], amt[3], tmp_4[12]);
	my_mux my_mux117(tmp_3[11], tmp_3[3], amt[3], tmp_4[11]);
	my_mux my_mux118(tmp_3[10], tmp_3[2], amt[3], tmp_4[10]);
	my_mux my_mux119(tmp_3[9], tmp_3[1], amt[3], tmp_4[9]);
	my_mux my_mux120(tmp_3[8], tmp_3[0], amt[3], tmp_4[8]);
	my_mux my_mux121(tmp_3[7], zero, amt[3], tmp_4[7]);
	my_mux my_mux122(tmp_3[6], zero, amt[3], tmp_4[6]);
	my_mux my_mux123(tmp_3[5], zero, amt[3], tmp_4[5]);
	my_mux my_mux124(tmp_3[4], zero, amt[3], tmp_4[4]);
	my_mux my_mux125(tmp_3[3], zero, amt[3], tmp_4[3]);
	my_mux my_mux126(tmp_3[2], zero, amt[3], tmp_4[2]);
	my_mux my_mux127(tmp_3[1], zero, amt[3], tmp_4[1]);
	my_mux my_mux128(tmp_3[0], zero, amt[3], tmp_4[0]);
	
	// layer 5
	my_mux my_mux129(tmp_4[31], tmp_4[15], amt[4], cout[31]);
	my_mux my_mux130(tmp_4[30], tmp_4[14], amt[4], cout[30]);
	my_mux my_mux131(tmp_4[29], tmp_4[13], amt[4], cout[29]);
	my_mux my_mux132(tmp_4[28], tmp_4[12], amt[4], cout[28]);
	my_mux my_mux133(tmp_4[27], tmp_4[11], amt[4], cout[27]);
	my_mux my_mux134(tmp_4[26], tmp_4[10], amt[4], cout[26]);
	my_mux my_mux135(tmp_4[25], tmp_4[9], amt[4], cout[25]);
	my_mux my_mux136(tmp_4[24], tmp_4[8], amt[4], cout[24]);
	my_mux my_mux137(tmp_4[23], tmp_4[7], amt[4], cout[23]);
	my_mux my_mux138(tmp_4[22], tmp_4[6], amt[4], cout[22]);
	my_mux my_mux139(tmp_4[21], tmp_4[5], amt[4], cout[21]);
	my_mux my_mux140(tmp_4[20], tmp_4[4], amt[4], cout[20]);
	my_mux my_mux141(tmp_4[19], tmp_4[3], amt[4], cout[19]);
	my_mux my_mux142(tmp_4[18], tmp_4[2], amt[4], cout[18]);
	my_mux my_mux143(tmp_4[17], tmp_4[1], amt[4], cout[17]);
	my_mux my_mux144(tmp_4[16], tmp_4[0], amt[4], cout[16]);
	my_mux my_mux145(tmp_4[15], zero, amt[4], cout[15]);
	my_mux my_mux146(tmp_4[14], zero, amt[4], cout[14]);
	my_mux my_mux147(tmp_4[13], zero, amt[4], cout[13]);
	my_mux my_mux148(tmp_4[12], zero, amt[4], cout[12]);
	my_mux my_mux149(tmp_4[11], zero, amt[4], cout[11]);
	my_mux my_mux150(tmp_4[10], zero, amt[4], cout[10]);
	my_mux my_mux151(tmp_4[9], zero, amt[4], cout[9]);
	my_mux my_mux152(tmp_4[8], zero, amt[4], cout[8]);
	my_mux my_mux153(tmp_4[7], zero, amt[4], cout[7]);
	my_mux my_mux154(tmp_4[6], zero, amt[4], cout[6]);
	my_mux my_mux155(tmp_4[5], zero, amt[4], cout[5]);
	my_mux my_mux156(tmp_4[4], zero, amt[4], cout[4]);
	my_mux my_mux157(tmp_4[3], zero, amt[4], cout[3]);
	my_mux my_mux158(tmp_4[2], zero, amt[4], cout[2]);
	my_mux my_mux159(tmp_4[1], zero, amt[4], cout[1]);
	my_mux my_mux160(tmp_4[0], zero, amt[4], cout[0]);
	
endmodule