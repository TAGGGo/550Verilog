module my_not(a, cout);
	 input [31:0] a;
	 output [31:0] cout;
	 not mynot_0(cout[0], a[0]);
    not mynot_1(cout[1], a[1]);
    not mynot_2(cout[2], a[2]);
    not mynot_3(cout[3], a[3]);
    not mynot_4(cout[4], a[4]);
    not mynot_5(cout[5], a[5]);
    not mynot_6(cout[6], a[6]);
    not mynot_7(cout[7], a[7]);
    not mynot_8(cout[8], a[8]);
    not mynot_9(cout[9], a[9]);
    not mynot_10(cout[10], a[10]);
    not mynot_11(cout[11], a[11]);
    not mynot_12(cout[12], a[12]);
    not mynot_13(cout[13], a[13]);
    not mynot_14(cout[14], a[14]);
    not mynot_15(cout[15], a[15]);
    not mynot_16(cout[16], a[16]);
    not mynot_17(cout[17], a[17]);
    not mynot_18(cout[18], a[18]);
    not mynot_19(cout[19], a[19]);
    not mynot_20(cout[20], a[20]);
    not mynot_21(cout[21], a[21]);
    not mynot_22(cout[22], a[22]);
    not mynot_23(cout[23], a[23]);
    not mynot_24(cout[24], a[24]);
    not mynot_25(cout[25], a[25]);
    not mynot_26(cout[26], a[26]);
    not mynot_27(cout[27], a[27]);
    not mynot_28(cout[28], a[28]);
    not mynot_29(cout[29], a[29]);
    not mynot_30(cout[30], a[30]);
	 not mynot_31(cout[31], a[31]);
endmodule