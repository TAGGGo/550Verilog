module my_or(opA, opB, cout);
	input [31:0] opA, opB;
	output [31:0] cout;
	or my_or0(cout[0], opA[0], opB[0]);
	or my_or1(cout[1], opA[1], opB[1]);
	or my_or2(cout[2], opA[2], opB[2]);
	or my_or3(cout[3], opA[3], opB[3]);
	or my_or4(cout[4], opA[4], opB[4]);
	or my_or5(cout[5], opA[5], opB[5]);
	or my_or6(cout[6], opA[6], opB[6]);
	or my_or7(cout[7], opA[7], opB[7]);
	or my_or8(cout[8], opA[8], opB[8]);
	or my_or9(cout[9], opA[9], opB[9]);
	or my_or10(cout[10], opA[10], opB[10]);
	or my_or11(cout[11], opA[11], opB[11]);
	or my_or12(cout[12], opA[12], opB[12]);
	or my_or13(cout[13], opA[13], opB[13]);
	or my_or14(cout[14], opA[14], opB[14]);
	or my_or15(cout[15], opA[15], opB[15]);
	or my_or16(cout[16], opA[16], opB[16]);
	or my_or17(cout[17], opA[17], opB[17]);
	or my_or18(cout[18], opA[18], opB[18]);
	or my_or19(cout[19], opA[19], opB[19]);
	or my_or20(cout[20], opA[20], opB[20]);
	or my_or21(cout[21], opA[21], opB[21]);
	or my_or22(cout[22], opA[22], opB[22]);
	or my_or23(cout[23], opA[23], opB[23]);
	or my_or24(cout[24], opA[24], opB[24]);
	or my_or25(cout[25], opA[25], opB[25]);
	or my_or26(cout[26], opA[26], opB[26]);
	or my_or27(cout[27], opA[27], opB[27]);
	or my_or28(cout[28], opA[28], opB[28]);
	or my_or29(cout[29], opA[29], opB[29]);
	or my_or30(cout[30], opA[30], opB[30]);
	or my_or31(cout[31], opA[31], opB[31]);
endmodule